`timescale 1ns/1ps

module nmcu_tb;



endmodule